`timescale 1ns / 1ps

module Top(
    input clk,
    input rst
);

    // autowire required

endmodule // Top
