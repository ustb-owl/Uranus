`timescale 1ns / 1ps

module GPIO(
    input clk,
    input rst,
    // IO
    input en,
    input write_en,
);

endmodule // GPIO
