`timescale 1ns / 1ps

module Top(
    input clk,
    input rst,
    //
);

//

endmodule // Top
