`timescale 1ns / 1ps

module Uranus(
    input clk,
    input rst
);

    //

endmodule // Uranus
