`timescale 1ns / 1ps

module PC(
    input clk,
    input rst,
);

endmodule // PC