`timescale 1ns / 1ps

module TLB(
    input clk,
    input rst
);

endmodule // TLB
