`timescale 1ns / 1ps

module ROM(
    input en,
    input 
);

endmodule // ROM
